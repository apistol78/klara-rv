module CPU_PreDecode (
	i_reset,
	i_clock,
	i_data,
	o_data
);
	input i_reset;
	input i_clock;
	input wire [120:0] i_data;
	output wire [120:0] o_data;
	reg [120:0] data = 0;
	assign o_data = data;
	wire is_ADD = (i_data[119:88] & 32'hfe00707f) == 32'h00000033;
	wire is_ADDI = (i_data[103:88] & 16'h707f) == 16'h0013;
	wire is_AND = (i_data[119:88] & 32'hfe00707f) == 32'h00007033;
	wire is_ANDI = (i_data[103:88] & 16'h707f) == 16'h7013;
	wire is_AUIPC = (i_data[95:88] & 8'h7f) == 8'h17;
	wire is_BEQ = (i_data[103:88] & 16'h707f) == 16'h0063;
	wire is_BGE = (i_data[103:88] & 16'h707f) == 16'h5063;
	wire is_BGEU = (i_data[103:88] & 16'h707f) == 16'h7063;
	wire is_BLT = (i_data[103:88] & 16'h707f) == 16'h4063;
	wire is_BLTU = (i_data[103:88] & 16'h707f) == 16'h6063;
	wire is_BNE = (i_data[103:88] & 16'h707f) == 16'h1063;
	wire is_CSRRC = (i_data[103:88] & 16'h707f) == 16'h3073;
	wire is_CSRRS = (i_data[103:88] & 16'h707f) == 16'h2073;
	wire is_CSRRW = (i_data[103:88] & 16'h707f) == 16'h1073;
	wire is_DIV = (i_data[119:88] & 32'hfe00707f) == 32'h02004033;
	wire is_DIVU = (i_data[119:88] & 32'hfe00707f) == 32'h02005033;
	wire is_EBREAK = (i_data[119:88] & 32'hffffffff) == 32'h00100073;
	wire is_ECALL = (i_data[119:88] & 32'hffffffff) == 32'h00000073;
	wire is_FADD = (i_data[119:88] & 32'hfe00007f) == 32'h00000053;
	wire is_FCVT_W_S = (i_data[119:88] & 32'hfff0007f) == 32'hc0000053;
	wire is_FCVT_WU_S = (i_data[119:88] & 32'hfff0007f) == 32'hc0100053;
	wire is_FCVT_S_W = (i_data[119:88] & 32'hfff0007f) == 32'hd0000053;
	wire is_FCVT_S_WU = (i_data[119:88] & 32'hfff0007f) == 32'hd0100053;
	wire is_FDIV = (i_data[119:88] & 32'hfe00007f) == 32'h18000053;
	wire is_FENCE = (i_data[103:88] & 16'h707f) == 16'h000f;
	wire is_FEQ = (i_data[119:88] & 32'hfe00707f) == 32'ha0002053;
	wire is_FLE = (i_data[119:88] & 32'hfe00707f) == 32'ha0000053;
	wire is_FLT = (i_data[119:88] & 32'hfe00707f) == 32'ha0001053;
	wire is_FLW = (i_data[103:88] & 16'h707f) == 16'h2007;
	wire is_FMADD = (i_data[119:88] & 32'h0600007f) == 32'h00000043;
	wire is_FMSUB = (i_data[119:88] & 32'h0600007f) == 32'h00000047;
	wire is_FNMADD = (i_data[119:88] & 32'h0600007f) == 32'h0000004f;
	wire is_FNMSUB = (i_data[119:88] & 32'h0600007f) == 32'h0000004b;
	wire is_FMIN = (i_data[119:88] & 32'hfe00707f) == 32'h28000053;
	wire is_FMAX = (i_data[119:88] & 32'hfe00707f) == 32'h28001053;
	wire is_FMUL = (i_data[119:88] & 32'hfe00007f) == 32'h10000053;
	wire is_FMV_X_W = (i_data[119:88] & 32'hfff0707f) == 32'he0000053;
	wire is_FMV_W_X = (i_data[119:88] & 32'hfff0707f) == 32'hf0000053;
	wire is_FSGNJ = (i_data[119:88] & 32'hfe00707f) == 32'h20000053;
	wire is_FSGNJN = (i_data[119:88] & 32'hfe00707f) == 32'h20001053;
	wire is_FSGNJX = (i_data[119:88] & 32'hfe00707f) == 32'h20002053;
	wire is_FSUB = (i_data[119:88] & 32'hfe00007f) == 32'h08000053;
	wire is_FSW = (i_data[103:88] & 16'h707f) == 16'h2027;
	wire is_JAL = (i_data[95:88] & 8'h7f) == 8'h6f;
	wire is_JALR = (i_data[103:88] & 16'h707f) == 16'h0067;
	wire is_LB = (i_data[103:88] & 16'h707f) == 16'h0003;
	wire is_LBU = (i_data[103:88] & 16'h707f) == 16'h4003;
	wire is_LH = (i_data[103:88] & 16'h707f) == 16'h1003;
	wire is_LHU = (i_data[103:88] & 16'h707f) == 16'h5003;
	wire is_LUI = (i_data[95:88] & 8'h7f) == 8'h37;
	wire is_LW = (i_data[103:88] & 16'h707f) == 16'h2003;
	wire is_MUL = (i_data[119:88] & 32'hfe00707f) == 32'h02000033;
	wire is_MULH = (i_data[119:88] & 32'hfe00707f) == 32'h02001033;
	wire is_MULHU = (i_data[119:88] & 32'hfe00707f) == 32'h02003033;
	wire is_MRET = (i_data[119:88] & 32'hffffffff) == 32'h30200073;
	wire is_OR = (i_data[119:88] & 32'hfe00707f) == 32'h00006033;
	wire is_ORI = (i_data[103:88] & 16'h707f) == 16'h6013;
	wire is_REM = (i_data[119:88] & 32'hfe00707f) == 32'h02006033;
	wire is_REMU = (i_data[119:88] & 32'hfe00707f) == 32'h02007033;
	wire is_SB = (i_data[103:88] & 16'h707f) == 16'h0023;
	wire is_SH = (i_data[103:88] & 16'h707f) == 16'h1023;
	wire is_SLL = (i_data[119:88] & 32'hfe00707f) == 32'h00001033;
	wire is_SLLI = (i_data[119:88] & 32'hfc00707f) == 32'h00001013;
	wire is_SLT = (i_data[119:88] & 32'hfe00707f) == 32'h00002033;
	wire is_SLTI = (i_data[103:88] & 16'h707f) == 16'h2013;
	wire is_SLTIU = (i_data[103:88] & 16'h707f) == 16'h3013;
	wire is_SLTU = (i_data[119:88] & 32'hfe00707f) == 32'h00003033;
	wire is_SRA = (i_data[119:88] & 32'hfe00707f) == 32'h40005033;
	wire is_SRAI = (i_data[119:88] & 32'hfc00707f) == 32'h40005013;
	wire is_SRL = (i_data[119:88] & 32'hfe00707f) == 32'h00005033;
	wire is_SRLI = (i_data[119:88] & 32'hfc00707f) == 32'h00005013;
	wire is_SUB = (i_data[119:88] & 32'hfe00707f) == 32'h40000033;
	wire is_SW = (i_data[103:88] & 16'h707f) == 16'h2023;
	wire is_WFI = (i_data[119:88] & 32'hffffffff) == 32'h10500073;
	wire is_XOR = (i_data[119:88] & 32'hfe00707f) == 32'h00004033;
	wire is_XORI = (i_data[103:88] & 16'h707f) == 16'h4013;
	wire is_B = ((((is_BEQ | is_BGE) | is_BGEU) | is_BLT) | is_BLTU) | is_BNE;
	wire is_I = ((((((((((((is_ADDI | is_ANDI) | is_FENCE) | is_FLW) | is_JALR) | is_LB) | is_LBU) | is_LH) | is_LHU) | is_LW) | is_ORI) | is_SLTI) | is_SLTIU) | is_XORI;
	wire is_J = is_JAL;
	wire is_R = ((((((((((((((((((((((((((((((((((((is_ADD | is_AND) | is_DIV) | is_DIVU) | is_FADD) | is_FCVT_W_S) | is_FCVT_WU_S) | is_FCVT_S_W) | is_FCVT_S_WU) | is_FDIV) | is_FEQ) | is_FLE) | is_FLT) | is_FMIN) | is_FMAX) | is_FMUL) | is_FMV_X_W) | is_FMV_W_X) | is_FSGNJ) | is_FSGNJN) | is_FSGNJX) | is_FSUB) | is_MUL) | is_MULH) | is_MULHU) | is_OR) | is_REM) | is_REMU) | is_SLL) | is_SLLI) | is_SLT) | is_SLTU) | is_SRA) | is_SRAI) | is_SRL) | is_SRLI) | is_SUB) | is_XOR;
	wire is_R4 = ((is_FMADD | is_FMSUB) | is_FNMADD) | is_FNMSUB;
	wire is_S = ((is_FSW | is_SB) | is_SH) | is_SW;
	wire is_U = is_AUIPC | is_LUI;
	wire is_CSR = ((is_CSRRC | is_CSRRS) | is_CSRRW) | is_MRET;
	wire is_ARITHMETIC = (((((((((is_ADD | is_ADDI) | is_AND) | is_ANDI) | is_AUIPC) | is_LUI) | is_OR) | is_ORI) | is_SUB) | is_XOR) | is_XORI;
	wire is_SHIFT = ((((is_SLL | is_SLLI) | is_SRA) | is_SRAI) | is_SRL) | is_SRLI;
	wire is_COMPARE = ((is_SLT | is_SLTI) | is_SLTIU) | is_SLTU;
	wire is_COMPLEX = (((((((((((((is_CSRRC | is_CSRRS) | is_CSRRW) | is_DIV) | is_DIVU) | is_EBREAK) | is_ECALL) | is_FENCE) | is_MUL) | is_MULH) | is_MULHU) | is_MRET) | is_REM) | is_REMU) | is_WFI;
	wire is_JUMP = is_JAL | is_JALR;
	wire is_JUMP_CONDITIONAL = ((((is_BEQ | is_BGE) | is_BGEU) | is_BLT) | is_BLTU) | is_BNE;
	wire is_MEMORY = ((((((is_LB | is_LBU) | is_LH) | is_LHU) | is_LW) | is_SB) | is_SH) | is_SW;
	wire is_FPU = ((((((((((((((((((((is_FADD | is_FCVT_W_S) | is_FCVT_WU_S) | is_FCVT_S_W) | is_FCVT_S_WU) | is_FDIV) | is_FEQ) | is_FLE) | is_FLT) | is_FMADD) | is_FMSUB) | is_FNMADD) | is_FNMSUB) | is_FMIN) | is_FMAX) | is_FMUL) | is_FMV_X_W) | is_FMV_W_X) | is_FSGNJ) | is_FSGNJN) | is_FSGNJX) | is_FSUB;
	wire is_FPU_MEMORY = is_FLW | is_FSW;
	wire RD_bank = (is_FADD ? 1'd1 : (is_FCVT_S_W ? 1'd1 : (is_FCVT_S_WU ? 1'd1 : (is_FDIV ? 1'd1 : (is_FLW ? 1'd1 : (is_FMADD ? 1'd1 : (is_FMSUB ? 1'd1 : (is_FNMADD ? 1'd1 : (is_FNMSUB ? 1'd1 : (is_FMIN ? 1'd1 : (is_FMAX ? 1'd1 : (is_FMUL ? 1'd1 : (is_FMV_W_X ? 1'd1 : (is_FSGNJ ? 1'd1 : (is_FSGNJN ? 1'd1 : (is_FSGNJX ? 1'd1 : (is_FSUB ? 1'd1 : 1'b0)))))))))))))))));
	wire RS1_bank = (is_FADD ? 1'd1 : (is_FCVT_W_S ? 1'd1 : (is_FCVT_WU_S ? 1'd1 : (is_FDIV ? 1'd1 : (is_FEQ ? 1'd1 : (is_FLE ? 1'd1 : (is_FLT ? 1'd1 : (is_FMADD ? 1'd1 : (is_FMSUB ? 1'd1 : (is_FNMADD ? 1'd1 : (is_FNMSUB ? 1'd1 : (is_FMIN ? 1'd1 : (is_FMAX ? 1'd1 : (is_FMUL ? 1'd1 : (is_FMV_X_W ? 1'd1 : (is_FSGNJ ? 1'd1 : (is_FSGNJN ? 1'd1 : (is_FSGNJX ? 1'd1 : (is_FSUB ? 1'd1 : 1'b0)))))))))))))))))));
	wire RS2_bank = (is_FADD ? 1'd1 : (is_FDIV ? 1'd1 : (is_FEQ ? 1'd1 : (is_FLE ? 1'd1 : (is_FLT ? 1'd1 : (is_FMADD ? 1'd1 : (is_FMSUB ? 1'd1 : (is_FNMADD ? 1'd1 : (is_FNMSUB ? 1'd1 : (is_FMIN ? 1'd1 : (is_FMAX ? 1'd1 : (is_FMUL ? 1'd1 : (is_FSGNJ ? 1'd1 : (is_FSGNJN ? 1'd1 : (is_FSGNJX ? 1'd1 : (is_FSUB ? 1'd1 : (is_FSW ? 1'd1 : 1'b0)))))))))))))))));
	wire RS3_bank = (is_FMADD ? 1'd1 : (is_FMSUB ? 1'd1 : (is_FNMADD ? 1'd1 : (is_FNMSUB ? 1'd1 : 1'b0))));
	wire have_RS1 = ((((is_B | is_I) | is_R) | is_S) | is_CSR) | is_R4;
	wire have_RS2 = ((is_B | is_R) | is_S) | is_R4;
	wire have_RS3 = is_R4;
	wire have_RD = ((((is_I | is_J) | is_R) | is_U) | is_CSR) | is_R4;
	wire [31:0] inst_B_imm = {{20 {i_data[119]}}, i_data[95], i_data[118:113], i_data[99:96], 1'b0};
	wire [31:0] inst_I_imm = {{21 {i_data[119]}}, i_data[118:108]};
	wire [31:0] inst_J_imm = {{12 {i_data[119]}}, i_data[107:100], i_data[108], i_data[118:109], 1'b0};
	wire [31:0] inst_S_imm = {{21 {i_data[119]}}, i_data[118:113], i_data[99:95]};
	wire [31:0] inst_U_imm = {i_data[119:100], 12'b000000000000};
	wire [31:0] inst_R_imm = {26'b00000000000000000000000000, i_data[113:108]};
	wire [31:0] inst_CSR_imm = {20'b00000000000000000000, i_data[119:108]};
	function automatic [5:0] sv2v_cast_6;
		input reg [5:0] inp;
		sv2v_cast_6 = inp;
	endfunction
	always @(posedge i_clock)
		if (i_reset)
			data <= 0;
		else begin
			data <= i_data;
			data[55-:6] <= sv2v_cast_6((have_RS1 ? {i_data[107:103]} : 5'h00));
			data[49-:6] <= sv2v_cast_6((have_RS2 ? {i_data[112:108]} : 5'h00));
			data[37-:6] <= sv2v_cast_6((have_RD ? {i_data[99:95]} : 5'h00));
			data[31-:32] <= (is_B ? inst_B_imm : (is_I ? inst_I_imm : (is_J ? inst_J_imm : (is_S ? inst_S_imm : (is_U ? inst_U_imm : (is_R ? inst_R_imm : (is_CSR ? inst_CSR_imm : 32'h00000000)))))));
		end
endmodule