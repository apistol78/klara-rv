module CPU_Decode (
	i_reset,
	i_clock,
	o_fault,
	i_data,
	o_data
);
	input i_reset;
	input i_clock;
	output reg o_fault;
	input wire [120:0] i_data;
	output wire [127:0] o_data;
	localparam OP_CSRRC = 4'd1;
	localparam OP_CSRRS = 4'd2;
	localparam OP_CSRRW = 4'd3;
	localparam OP_DIV = 4'd4;
	localparam OP_DIVU = 4'd5;
	localparam OP_EBREAK = 4'd6;
	localparam OP_ECALL = 4'd7;
	localparam OP_FENCE = 4'd8;
	localparam OP_MUL = 4'd9;
	localparam OP_MULH = 4'd10;
	localparam OP_MULHU = 4'd11;
	localparam OP_MRET = 4'd12;
	localparam OP_REM = 4'd13;
	localparam OP_REMU = 4'd14;
	wire is_ADD = (i_data[119:88] & 32'hfe00707f) == 32'h00000033;
	wire is_ADDI = (i_data[103:88] & 16'h707f) == 16'h0013;
	wire is_AND = (i_data[119:88] & 32'hfe00707f) == 32'h00007033;
	wire is_ANDI = (i_data[103:88] & 16'h707f) == 16'h7013;
	wire is_AUIPC = (i_data[95:88] & 8'h7f) == 8'h17;
	wire is_BEQ = (i_data[103:88] & 16'h707f) == 16'h0063;
	wire is_BGE = (i_data[103:88] & 16'h707f) == 16'h5063;
	wire is_BGEU = (i_data[103:88] & 16'h707f) == 16'h7063;
	wire is_BLT = (i_data[103:88] & 16'h707f) == 16'h4063;
	wire is_BLTU = (i_data[103:88] & 16'h707f) == 16'h6063;
	wire is_BNE = (i_data[103:88] & 16'h707f) == 16'h1063;
	wire is_CSRRC = (i_data[103:88] & 16'h707f) == 16'h3073;
	wire is_CSRRS = (i_data[103:88] & 16'h707f) == 16'h2073;
	wire is_CSRRW = (i_data[103:88] & 16'h707f) == 16'h1073;
	wire is_DIV = (i_data[119:88] & 32'hfe00707f) == 32'h02004033;
	wire is_DIVU = (i_data[119:88] & 32'hfe00707f) == 32'h02005033;
	wire is_EBREAK = (i_data[119:88] & 32'hffffffff) == 32'h00100073;
	wire is_ECALL = (i_data[119:88] & 32'hffffffff) == 32'h00000073;
	wire is_FADD = (i_data[119:88] & 32'hfe00007f) == 32'h00000053;
	wire is_FCVT_W_S = (i_data[119:88] & 32'hfff0007f) == 32'hc0000053;
	wire is_FCVT_WU_S = (i_data[119:88] & 32'hfff0007f) == 32'hc0100053;
	wire is_FCVT_S_W = (i_data[119:88] & 32'hfff0007f) == 32'hd0000053;
	wire is_FCVT_S_WU = (i_data[119:88] & 32'hfff0007f) == 32'hd0100053;
	wire is_FDIV = (i_data[119:88] & 32'hfe00007f) == 32'h18000053;
	wire is_FENCE = (i_data[103:88] & 16'h707f) == 16'h000f;
	wire is_FEQ = (i_data[119:88] & 32'hfe00707f) == 32'ha0002053;
	wire is_FLE = (i_data[119:88] & 32'hfe00707f) == 32'ha0000053;
	wire is_FLT = (i_data[119:88] & 32'hfe00707f) == 32'ha0001053;
	wire is_FLW = (i_data[103:88] & 16'h707f) == 16'h2007;
	wire is_FMADD = (i_data[119:88] & 32'h0600007f) == 32'h00000043;
	wire is_FMSUB = (i_data[119:88] & 32'h0600007f) == 32'h00000047;
	wire is_FNMADD = (i_data[119:88] & 32'h0600007f) == 32'h0000004f;
	wire is_FNMSUB = (i_data[119:88] & 32'h0600007f) == 32'h0000004b;
	wire is_FMIN = (i_data[119:88] & 32'hfe00707f) == 32'h28000053;
	wire is_FMAX = (i_data[119:88] & 32'hfe00707f) == 32'h28001053;
	wire is_FMUL = (i_data[119:88] & 32'hfe00007f) == 32'h10000053;
	wire is_FMV_X_W = (i_data[119:88] & 32'hfff0707f) == 32'he0000053;
	wire is_FMV_W_X = (i_data[119:88] & 32'hfff0707f) == 32'hf0000053;
	wire is_FSGNJ = (i_data[119:88] & 32'hfe00707f) == 32'h20000053;
	wire is_FSGNJN = (i_data[119:88] & 32'hfe00707f) == 32'h20001053;
	wire is_FSGNJX = (i_data[119:88] & 32'hfe00707f) == 32'h20002053;
	wire is_FSUB = (i_data[119:88] & 32'hfe00007f) == 32'h08000053;
	wire is_FSW = (i_data[103:88] & 16'h707f) == 16'h2027;
	wire is_JAL = (i_data[95:88] & 8'h7f) == 8'h6f;
	wire is_JALR = (i_data[103:88] & 16'h707f) == 16'h0067;
	wire is_LB = (i_data[103:88] & 16'h707f) == 16'h0003;
	wire is_LBU = (i_data[103:88] & 16'h707f) == 16'h4003;
	wire is_LH = (i_data[103:88] & 16'h707f) == 16'h1003;
	wire is_LHU = (i_data[103:88] & 16'h707f) == 16'h5003;
	wire is_LUI = (i_data[95:88] & 8'h7f) == 8'h37;
	wire is_LW = (i_data[103:88] & 16'h707f) == 16'h2003;
	wire is_MUL = (i_data[119:88] & 32'hfe00707f) == 32'h02000033;
	wire is_MULH = (i_data[119:88] & 32'hfe00707f) == 32'h02001033;
	wire is_MULHU = (i_data[119:88] & 32'hfe00707f) == 32'h02003033;
	wire is_MRET = (i_data[119:88] & 32'hffffffff) == 32'h30200073;
	wire is_OR = (i_data[119:88] & 32'hfe00707f) == 32'h00006033;
	wire is_ORI = (i_data[103:88] & 16'h707f) == 16'h6013;
	wire is_REM = (i_data[119:88] & 32'hfe00707f) == 32'h02006033;
	wire is_REMU = (i_data[119:88] & 32'hfe00707f) == 32'h02007033;
	wire is_SB = (i_data[103:88] & 16'h707f) == 16'h0023;
	wire is_SH = (i_data[103:88] & 16'h707f) == 16'h1023;
	wire is_SLL = (i_data[119:88] & 32'hfe00707f) == 32'h00001033;
	wire is_SLLI = (i_data[119:88] & 32'hfc00707f) == 32'h00001013;
	wire is_SLT = (i_data[119:88] & 32'hfe00707f) == 32'h00002033;
	wire is_SLTI = (i_data[103:88] & 16'h707f) == 16'h2013;
	wire is_SLTIU = (i_data[103:88] & 16'h707f) == 16'h3013;
	wire is_SLTU = (i_data[119:88] & 32'hfe00707f) == 32'h00003033;
	wire is_SRA = (i_data[119:88] & 32'hfe00707f) == 32'h40005033;
	wire is_SRAI = (i_data[119:88] & 32'hfc00707f) == 32'h40005013;
	wire is_SRL = (i_data[119:88] & 32'hfe00707f) == 32'h00005033;
	wire is_SRLI = (i_data[119:88] & 32'hfc00707f) == 32'h00005013;
	wire is_SUB = (i_data[119:88] & 32'hfe00707f) == 32'h40000033;
	wire is_SW = (i_data[103:88] & 16'h707f) == 16'h2023;
	wire is_WFI = (i_data[119:88] & 32'hffffffff) == 32'h10500073;
	wire is_XOR = (i_data[119:88] & 32'hfe00707f) == 32'h00004033;
	wire is_XORI = (i_data[103:88] & 16'h707f) == 16'h4013;
	wire is_B = ((((is_BEQ | is_BGE) | is_BGEU) | is_BLT) | is_BLTU) | is_BNE;
	wire is_I = ((((((((((((is_ADDI | is_ANDI) | is_FENCE) | is_FLW) | is_JALR) | is_LB) | is_LBU) | is_LH) | is_LHU) | is_LW) | is_ORI) | is_SLTI) | is_SLTIU) | is_XORI;
	wire is_J = is_JAL;
	wire is_R = ((((((((((((((((((((((((((((((((((((is_ADD | is_AND) | is_DIV) | is_DIVU) | is_FADD) | is_FCVT_W_S) | is_FCVT_WU_S) | is_FCVT_S_W) | is_FCVT_S_WU) | is_FDIV) | is_FEQ) | is_FLE) | is_FLT) | is_FMIN) | is_FMAX) | is_FMUL) | is_FMV_X_W) | is_FMV_W_X) | is_FSGNJ) | is_FSGNJN) | is_FSGNJX) | is_FSUB) | is_MUL) | is_MULH) | is_MULHU) | is_OR) | is_REM) | is_REMU) | is_SLL) | is_SLLI) | is_SLT) | is_SLTU) | is_SRA) | is_SRAI) | is_SRL) | is_SRLI) | is_SUB) | is_XOR;
	wire is_R4 = ((is_FMADD | is_FMSUB) | is_FNMADD) | is_FNMSUB;
	wire is_S = ((is_FSW | is_SB) | is_SH) | is_SW;
	wire is_U = is_AUIPC | is_LUI;
	wire is_CSR = ((is_CSRRC | is_CSRRS) | is_CSRRW) | is_MRET;
	wire is_ARITHMETIC = (((((((((is_ADD | is_ADDI) | is_AND) | is_ANDI) | is_AUIPC) | is_LUI) | is_OR) | is_ORI) | is_SUB) | is_XOR) | is_XORI;
	wire is_SHIFT = ((((is_SLL | is_SLLI) | is_SRA) | is_SRAI) | is_SRL) | is_SRLI;
	wire is_COMPARE = ((is_SLT | is_SLTI) | is_SLTIU) | is_SLTU;
	wire is_COMPLEX = (((((((((((((is_CSRRC | is_CSRRS) | is_CSRRW) | is_DIV) | is_DIVU) | is_EBREAK) | is_ECALL) | is_FENCE) | is_MUL) | is_MULH) | is_MULHU) | is_MRET) | is_REM) | is_REMU) | is_WFI;
	wire is_JUMP = is_JAL | is_JALR;
	wire is_JUMP_CONDITIONAL = ((((is_BEQ | is_BGE) | is_BGEU) | is_BLT) | is_BLTU) | is_BNE;
	wire is_MEMORY = ((((((is_LB | is_LBU) | is_LH) | is_LHU) | is_LW) | is_SB) | is_SH) | is_SW;
	wire is_FPU = ((((((((((((((((((((is_FADD | is_FCVT_W_S) | is_FCVT_WU_S) | is_FCVT_S_W) | is_FCVT_S_WU) | is_FDIV) | is_FEQ) | is_FLE) | is_FLT) | is_FMADD) | is_FMSUB) | is_FNMADD) | is_FNMSUB) | is_FMIN) | is_FMAX) | is_FMUL) | is_FMV_X_W) | is_FMV_W_X) | is_FSGNJ) | is_FSGNJN) | is_FSGNJX) | is_FSUB;
	wire is_FPU_MEMORY = is_FLW | is_FSW;
	wire RD_bank = (is_FADD ? 1'd1 : (is_FCVT_S_W ? 1'd1 : (is_FCVT_S_WU ? 1'd1 : (is_FDIV ? 1'd1 : (is_FLW ? 1'd1 : (is_FMADD ? 1'd1 : (is_FMSUB ? 1'd1 : (is_FNMADD ? 1'd1 : (is_FNMSUB ? 1'd1 : (is_FMIN ? 1'd1 : (is_FMAX ? 1'd1 : (is_FMUL ? 1'd1 : (is_FMV_W_X ? 1'd1 : (is_FSGNJ ? 1'd1 : (is_FSGNJN ? 1'd1 : (is_FSGNJX ? 1'd1 : (is_FSUB ? 1'd1 : 1'b0)))))))))))))))));
	wire RS1_bank = (is_FADD ? 1'd1 : (is_FCVT_W_S ? 1'd1 : (is_FCVT_WU_S ? 1'd1 : (is_FDIV ? 1'd1 : (is_FEQ ? 1'd1 : (is_FLE ? 1'd1 : (is_FLT ? 1'd1 : (is_FMADD ? 1'd1 : (is_FMSUB ? 1'd1 : (is_FNMADD ? 1'd1 : (is_FNMSUB ? 1'd1 : (is_FMIN ? 1'd1 : (is_FMAX ? 1'd1 : (is_FMUL ? 1'd1 : (is_FMV_X_W ? 1'd1 : (is_FSGNJ ? 1'd1 : (is_FSGNJN ? 1'd1 : (is_FSGNJX ? 1'd1 : (is_FSUB ? 1'd1 : 1'b0)))))))))))))))))));
	wire RS2_bank = (is_FADD ? 1'd1 : (is_FDIV ? 1'd1 : (is_FEQ ? 1'd1 : (is_FLE ? 1'd1 : (is_FLT ? 1'd1 : (is_FMADD ? 1'd1 : (is_FMSUB ? 1'd1 : (is_FNMADD ? 1'd1 : (is_FNMSUB ? 1'd1 : (is_FMIN ? 1'd1 : (is_FMAX ? 1'd1 : (is_FMUL ? 1'd1 : (is_FSGNJ ? 1'd1 : (is_FSGNJN ? 1'd1 : (is_FSGNJX ? 1'd1 : (is_FSUB ? 1'd1 : (is_FSW ? 1'd1 : 1'b0)))))))))))))))));
	wire RS3_bank = (is_FMADD ? 1'd1 : (is_FMSUB ? 1'd1 : (is_FNMADD ? 1'd1 : (is_FNMSUB ? 1'd1 : 1'b0))));
	wire [3:0] alu_operation = (is_ADD ? 0 : (is_ADDI ? 0 : (is_AND ? 3 : (is_ANDI ? 3 : (is_AUIPC ? 0 : (is_BEQ ? 11 : (is_BGE ? 13 : (is_BGEU ? 14 : (is_BLT ? 9 : (is_BLTU ? 10 : (is_BNE ? 12 : (is_FLW ? 0 : (is_FSW ? 0 : (is_JAL ? 0 : (is_JALR ? 0 : (is_LB ? 0 : (is_LBU ? 0 : (is_LH ? 0 : (is_LHU ? 0 : (is_LUI ? 1 : (is_LW ? 0 : (is_OR ? 4 : (is_ORI ? 4 : (is_SB ? 0 : (is_SH ? 0 : (is_SLL ? 6 : (is_SLLI ? 6 : (is_SLT ? 9 : (is_SLTI ? 9 : (is_SLTIU ? 10 : (is_SLTU ? 10 : (is_SRA ? 8 : (is_SRAI ? 8 : (is_SRL ? 7 : (is_SRLI ? 7 : (is_SUB ? 2 : (is_SW ? 0 : (is_XOR ? 5 : (is_XORI ? 5 : 4'd0)))))))))))))))))))))))))))))))))))))));
	wire [4:0] alu_operand1 = (is_AUIPC ? 5'b01000 : (is_JAL ? 5'b01000 : (is_LUI ? 5'b10000 : 5'b00010)));
	wire [4:0] alu_operand2 = (is_ADDI ? 5'b10000 : (is_ANDI ? 5'b10000 : (is_AUIPC ? 5'b10000 : (is_FLW ? 5'b10000 : (is_FSW ? 5'b10000 : (is_JAL ? 5'b10000 : (is_JALR ? 5'b10000 : (is_LB ? 5'b10000 : (is_LBU ? 5'b10000 : (is_LH ? 5'b10000 : (is_LHU ? 5'b10000 : (is_LUI ? 5'b00001 : (is_LW ? 5'b10000 : (is_ORI ? 5'b10000 : (is_SB ? 5'b10000 : (is_SH ? 5'b10000 : (is_SLLI ? 5'b10000 : (is_SLTI ? 5'b10000 : (is_SLTIU ? 5'b10000 : (is_SRAI ? 5'b10000 : (is_SRLI ? 5'b10000 : (is_SW ? 5'b10000 : (is_XORI ? 5'b10000 : 5'b00100)))))))))))))))))))))));
	wire memory_read = (((((is_FLW | is_LB) | is_LBU) | is_LH) | is_LHU) | is_LW) | 1'b0;
	wire memory_write = (((is_FSW | is_SB) | is_SH) | is_SW) | 1'b0;
	wire [1:0] memory_width = (is_FLW ? 2'b10 : (is_FSW ? 2'b10 : (is_LB ? 2'b00 : (is_LBU ? 2'b00 : (is_LH ? 2'b01 : (is_LHU ? 2'b01 : (is_LW ? 2'b10 : (is_SB ? 2'b00 : (is_SH ? 2'b01 : (is_SW ? 2'b10 : 3'd0))))))))));
	wire memory_signed = (is_LB | is_LH) | 1'b0;
	wire [4:0] fpu_operation = (is_FADD ? 0 : (is_FCVT_W_S ? 8 : (is_FCVT_WU_S ? 9 : (is_FCVT_S_W ? 10 : (is_FCVT_S_WU ? 11 : (is_FDIV ? 3 : (is_FEQ ? 13 : (is_FLE ? 15 : (is_FLT ? 14 : (is_FMADD ? 4 : (is_FMSUB ? 5 : (is_FNMADD ? 6 : (is_FNMSUB ? 7 : (is_FMIN ? 19 : (is_FMAX ? 20 : (is_FMUL ? 2 : (is_FMV_X_W ? 12 : (is_FMV_W_X ? 12 : (is_FSGNJ ? 16 : (is_FSGNJN ? 17 : (is_FSGNJX ? 18 : (is_FSUB ? 1 : 5'd0))))))))))))))))))))));
	wire have_RS1 = ((((is_B | is_I) | is_R) | is_S) | is_CSR) | is_R4;
	wire have_RS2 = ((is_B | is_R) | is_S) | is_R4;
	wire have_RS3 = is_R4;
	wire have_RD = ((((is_I | is_J) | is_R) | is_U) | is_CSR) | is_R4;
	wire [31:0] inst_B_imm = {{20 {i_data[119]}}, i_data[95], i_data[118:113], i_data[99:96], 1'b0};
	wire [31:0] inst_I_imm = {{21 {i_data[119]}}, i_data[118:108]};
	wire [31:0] inst_J_imm = {{12 {i_data[119]}}, i_data[107:100], i_data[108], i_data[118:109], 1'b0};
	wire [31:0] inst_S_imm = {{21 {i_data[119]}}, i_data[118:113], i_data[99:95]};
	wire [31:0] inst_U_imm = {i_data[119:100], 12'b000000000000};
	wire [31:0] inst_R_imm = {26'b00000000000000000000000000, i_data[113:108]};
	wire [31:0] inst_CSR_imm = {20'b00000000000000000000, i_data[119:108]};
	reg [127:0] data = 0;
	assign o_data = data;
	initial o_fault = 0;
	always @(posedge i_clock)
		if (i_reset) begin
			data <= 0;
			o_fault <= 0;
		end
		else begin
			data[126-:32] <= i_data[87-:32];
			data[94-:3] <= {(i_data[43-:6] != 0 ? 1'b1 : 1'b0), (i_data[49-:6] != 0 ? 1'b1 : 1'b0), (i_data[55-:6] != 0 ? 1'b1 : 1'b0)};
			data[91-:6] <= i_data[55-:6];
			data[85-:6] <= i_data[49-:6];
			data[79-:6] <= i_data[43-:6];
			data[73-:6] <= i_data[37-:6];
			data[67-:32] <= (is_B ? inst_B_imm : (is_I ? inst_I_imm : (is_J ? inst_J_imm : (is_S ? inst_S_imm : (is_U ? inst_U_imm : (is_R ? inst_R_imm : (is_CSR ? inst_CSR_imm : 32'h00000000)))))));
			data[35] <= is_ARITHMETIC;
			data[34] <= is_SHIFT;
			data[33] <= is_COMPARE;
			data[32] <= is_COMPLEX;
			data[31] <= is_JUMP;
			data[30] <= is_JUMP_CONDITIONAL;
			data[29-:4] <= alu_operation;
			data[25-:5] <= alu_operand1;
			data[20-:5] <= alu_operand2;
			data[15] <= memory_read;
			data[14] <= memory_write;
			data[13-:2] <= memory_width;
			data[11] <= memory_signed;
			data[5] <= is_FPU;
			data[4-:5] <= fpu_operation;
			data[10-:5] <= (is_CSRRC ? OP_CSRRC : (is_CSRRS ? OP_CSRRS : (is_CSRRW ? OP_CSRRW : (is_DIV ? OP_DIV : (is_DIVU ? OP_DIVU : (is_EBREAK ? OP_EBREAK : (is_ECALL ? OP_ECALL : (is_FENCE ? OP_FENCE : (is_MUL ? OP_MUL : (is_MULH ? OP_MULH : (is_MULHU ? OP_MULHU : (is_MRET ? OP_MRET : (is_REM ? OP_REM : (is_REMU ? OP_REMU : 0))))))))))))));
			data[127] <= i_data[120];
		end
endmodule