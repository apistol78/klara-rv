/*
 Klara-RV
 Copyright (c) 2025 Anders Pistol.

 This Source Code Form is subject to the terms of the Mozilla Public
 License, v. 2.0. If a copy of the MPL was not distributed with this
 file, You can obtain one at https://mozilla.org/MPL/2.0/.
*/

`timescale 1ns/1ns
`define FREQUENCY 25000000

(* top *)
module SoC(
      input CLOCK_p,
      output LED_p,
	  output IO_p,
	  input UART_RX,
	  output UART_TX
);
	wire clock;
	wire reset = 1'b0;


	// current 1.04 MhZ signal at 125 MHz

	// 125 MHz
	PLL_ECP5 #(
		.CLKI_DIV(1),
		.CLKFB_DIV(5),
		.CLKOP_DIV(5),
		.CLKOP_CPHASE(0)
	) pll(
		.i_clk(CLOCK_p),
		.o_clk1(clock),
		.o_clk2(),
		.o_clk_locked()
	);


	//assign LED_p = cpu_dbus_request;
	assign IO_p = pin_value;


	bit pin_value = 1'b0;
	wire pin_select;
	bit pin_ready = 1'b0;

	always @(posedge clock) begin
		if (bus_request && pin_select) begin
			pin_value <= bus_wdata[0];
			pin_ready <= 1'b1;
		end
		else begin
			pin_ready <= 1'b0;
		end
	end


	//====================================================
	// ROM
	wire rom_select;
	wire [31:0] rom_address;
	wire [31:0] rom_rdata;
	wire rom_ready;

	SoC_BROM rom(
		.i_clock(clock),
		.i_request(bus_request && rom_select),
		.i_address(rom_address),
		.o_rdata(rom_rdata),
		.o_ready(rom_ready)
	);


	//====================================================
	// RAM
	wire ram_select;
	wire [31:0] ram_address;
	wire [31:0] ram_wdata;
	wire [31:0] ram_rdata;
	wire ram_ready;

	BRAM #(
		.SIZE(32'h400)
	) ram(
		.i_clock(clock),
		.i_request(bus_request && ram_select),
		.i_rw(bus_rw),
		.i_address(ram_address),
		.i_wdata(ram_wdata),
		.o_rdata(ram_rdata),
		.o_ready(ram_ready),
		.o_valid()
	);


	//====================================================
	// UART
	wire uart_select;
	wire [1:0] uart_address;
	wire [31:0] uart_wdata;
	wire [31:0] uart_rdata;
	wire uart_ready;

	UART #(
		.PRESCALE(`FREQUENCY / (9600 * 8)),
		.RX_FIFO_DEPTH(512)
	) uart(
		.i_reset(reset),
		.i_clock(clock),
		.i_request(bus_request && uart_select),
		.i_rw(bus_rw),
		.i_address(uart_address),
		.i_wdata(uart_wdata),
		.o_rdata(uart_rdata),
		.o_ready(uart_ready),
		.o_interrupt(),
		// ---
		.UART_RX(UART_RX),
		.UART_TX(UART_TX)
	);


	//====================================================
	// Chip select
	assign rom_select = bus_address[31:28] == 4'h0;
	assign rom_address = { 4'h0, bus_address[27:0] };

	assign ram_select = bus_address[31:28] == 4'h1;
	assign ram_address = { 4'h0, bus_address[27:0] };
	assign ram_wdata = bus_wdata;

	assign uart_select = bus_address[31:28] == 4'h3;
	assign uart_address = { 4'h0, bus_address[27:0] };
	assign uart_wdata = bus_wdata;

	assign pin_select = bus_address[31:28] == 4'h4;

	assign bus_rdata =
		rom_select		? rom_rdata		:
		ram_select		? ram_rdata		:
		uart_select		? uart_rdata	:
		32'h00000000;

	assign bus_ready =
		rom_select		? rom_ready		:
		ram_select		? ram_ready		:
		uart_select		? uart_ready	:
		pin_select		? pin_ready		:
		1'b0;


	//====================================================
	// CPU BusMux
	wire bus_rw;
	wire bus_request;
	wire bus_ready;
	wire [31:0] bus_address;
	wire [31:0] bus_rdata;
	wire [31:0] bus_wdata;

	CPU_BusMux #(
		.REGISTERED(1)
	) bus(
		.i_reset(reset),
		.i_clock(clock),

		.o_bus_rw(bus_rw),
		.o_bus_request(bus_request),
		.i_bus_ready(bus_ready),
		.o_bus_address(bus_address),
		.i_bus_rdata(bus_rdata),
		.o_bus_wdata(bus_wdata),

		.i_pa_request(cpu_ibus_request),
		.o_pa_ready(cpu_ibus_ready),
		.i_pa_address(cpu_ibus_address),
		.o_pa_rdata(cpu_ibus_rdata),

		.i_pb_rw(cpu_dbus_rw),
		.i_pb_request(cpu_dbus_request),
		.o_pb_ready(cpu_dbus_ready),
		.i_pb_address(cpu_dbus_address),
		.o_pb_rdata(cpu_dbus_rdata),
		.i_pb_wdata(cpu_dbus_wdata)
	);


	//====================================================
	// CPU
	wire cpu_ibus_request;
	wire cpu_ibus_ready;
	wire [31:0] cpu_ibus_address;
	wire [31:0] cpu_ibus_rdata;
	wire cpu_dbus_rw;
	wire cpu_dbus_request;
	wire cpu_dbus_ready;
	wire [31:0] cpu_dbus_address;
	wire [31:0] cpu_dbus_rdata;
	wire [31:0] cpu_dbus_wdata;
	wire cpu_fault;

	CPU #(
		.FREQUENCY(`FREQUENCY),
		.DCACHE_SIZE(0),
		.DCACHE_REGISTERED(1),
		.ICACHE_SIZE(1),
		.ICACHE_REGISTERED(1)		
	) cpu(
		.i_reset(reset),
		.i_clock(clock),

		// Control
		.i_timer_interrupt(1'b0),
		.i_external_interrupt(1'b0),

		// Instruction bus
		.o_ibus_request(cpu_ibus_request),
		.i_ibus_ready(cpu_ibus_ready),
		.o_ibus_address(cpu_ibus_address),
		.i_ibus_rdata(cpu_ibus_rdata),

		// Data bus
		.o_dbus_rw(cpu_dbus_rw),
		.o_dbus_request(cpu_dbus_request),
		.i_dbus_ready(cpu_dbus_ready),
		.o_dbus_address(cpu_dbus_address),
		.i_dbus_rdata(cpu_dbus_rdata),
		.o_dbus_wdata(cpu_dbus_wdata),

		// Debug
		.o_icache_hit(),
		.o_icache_miss(),
		.o_dcache_hit(),
		.o_dcache_miss(),
		.o_execute_busy(),
		.o_memory_busy(),
		.o_fault(cpu_fault)
	);

endmodule
