/*
 Klara-RV
 Copyright (c) 2025 Anders Pistol.

 This Source Code Form is subject to the terms of the Mozilla Public
 License, v. 2.0. If a copy of the MPL was not distributed with this
 file, You can obtain one at https://mozilla.org/MPL/2.0/.
*/
`include "CPU_Defines.sv"

`timescale 1ns/1ns
`default_nettype none

module CPU_ICache_None(
	input wire i_reset,
	input wire i_clock,
	
	input wire [31:0] i_input_pc,
	output bit [31:0] o_rdata,
	output bit o_ready,
	input wire i_stall,

	// Bus
	output bit o_bus_request,
	input wire i_bus_ready,
	output wire [31:0] o_bus_address,
	input wire [31:0] i_bus_rdata,

	// Debug
	output wire [31:0] o_hit,
	output wire [31:0] o_miss
);

	typedef enum bit [1:0]
	{
		IDLE		= 2'd0,
		READ_BUS	= 2'd1
	} state_t;

	state_t next = IDLE;
	state_t state = IDLE;

	// Debug, only for verilated.
	assign o_hit = 0;
	assign o_miss = 0;

	assign o_bus_address = i_input_pc;
	
	always_comb begin
		next = state;
	
		o_ready = 0;
		o_rdata = 32'h0;
		o_bus_request = 0;

		case (state)
			IDLE: begin
				if (!i_stall) begin
					o_bus_request = 1;
					next = READ_BUS;
				end
			end

			READ_BUS: begin
				o_bus_request = 1;
				if (i_bus_ready) begin
					o_ready = 1;
					o_rdata = i_bus_rdata;
					next = IDLE;
				end
			end
		endcase

		if (i_reset) begin
			next = IDLE;
		end
	end

endmodule
